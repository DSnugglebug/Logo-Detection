
library ieee;
use ieee.std_logic_1164.all;

entity simple_dual_port_ram_single_clock is

	generic 
	(
		DATA_WIDTH : natural;
		DATA_NUM : natural
	);

	port 
	(
		clk	: in std_logic;
		raddr	: in natural range 0 to DATA_NUM - 1;
		waddr	: in natural range 0 to DATA_NUM - 1;
		data	: in std_logic_vector((DATA_WIDTH-1) downto 0);
		we		: in std_logic := '1';
		q		: out std_logic_vector((DATA_WIDTH -1) downto 0)
	);

end simple_dual_port_ram_single_clock;

architecture rtl of simple_dual_port_ram_single_clock is

	-- Build a 2-D array type for the RAM
	subtype word_t is std_logic_vector((DATA_WIDTH-1) downto 0);
	type memory_t is array(DATA_NUM-1 downto 0) of word_t;

	-- Declare the RAM signal.	
	signal ram : memory_t;

begin

	process(clk)
	begin
	if(rising_edge(clk)) then 
		if(we = '1') then
			ram(waddr) <= data;
		end if;
 
		-- On a read during a write to the same address, the read will
		-- return the OLD data at the address
		q <= ram(raddr);
	end if;
	end process;

end rtl;
